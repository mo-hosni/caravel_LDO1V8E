** sch_path:
*+ /home/ahmedreda/Project/AR_BGR_with_Enable_line/schematic/fullldoEnBias/fullldoenbiasx.sch
.subckt EF_LDOR1V8E vdd vss vo en
*.PININFO vdd:B vss:B vo:O en:I
x1 vdd vss en vss vss vss vss vss vss vss vss vss vdd vss vss vss vss vss vss o1 o2 vo
+ fullldoEn3p3_v1
x2 vdd o2 o1 vss sbcx3
.ends

* expanding   symbol:  Project/AR_BGR_with_Enable_line/schematic/fullldoEn/fullldoEn3p3_v1.sym # of
*+ pins=7
** sym_path: /home/ahmedreda/Project/AR_BGR_with_Enable_line/schematic/fullldoEn/fullldoEn3p3_v1.sym
** sch_path: /home/ahmedreda/Project/AR_BGR_with_Enable_line/schematic/fullldoEn/fullldoEn3p3_v1.sch
.subckt fullldoEn3p3_v1 vdd vss en trim[15] trim[14] trim[13] trim[12] trim[11] trim[10] trim[9]
+ trim[8] trim[7] trim[6] trim[5] trim[4] trim[3] trim[2] trim[1] trim[0] biasbgr biasldo vo
*.PININFO vdd:B vss:B en:I trim[15:0]:I vo:O biasbgr:O biasldo:O
x1 trim[15] trim[14] trim[13] trim[12] trim[11] trim[10] trim[9] trim[8] trim[7] trim[6] trim[5]
+ trim[4] trim[3] trim[2] trim[1] trim[0] vss biasbgr vdd biasldo vg vo fullldoxc_v2_1
x2 vdd en vg vss tg1x
.ends


* expanding   symbol:  Project/AR_BGR_with_Enable_line/schematic/bias-circuit/sbcx3.sym # of pins=4
** sym_path: /home/ahmedreda/Project/AR_BGR_with_Enable_line/schematic/bias-circuit/sbcx3.sym
** sch_path: /home/ahmedreda/Project/AR_BGR_with_Enable_line/schematic/bias-circuit/sbcx3.sch
.subckt sbcx3 vdd o2 o1 vss
*.PININFO vdd:B o1:O o2:O vss:B
XM12 vssup or vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=6 nf=1 m=2
XM1 or or vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=6 nf=1 m=2
XM11 o1 or vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=6 nf=1 m=2
XM14 o2 or vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=6 nf=1 m=2
XM7 vdd vdd vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=6 nf=1 m=4
XM19 vssup vssup vss vss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=6 nf=1 m=2
XM2 or vssup net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=6 nf=1 m=8
XM9 or or or vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=6 nf=1 m=4
XM8 vss vss vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=6 nf=1 m=4
XR7 vss net1 vss sky130_fd_pr__res_xhigh_po W=0.69  L=4 mult=1 m=1
XR1 vss vss vss sky130_fd_pr__res_xhigh_po W=0.69  L=4 mult=1 m=1
XR2 vss vss vss sky130_fd_pr__res_xhigh_po W=0.69  L=4 mult=1 m=1
XR3 net2 vdd vss sky130_fd_pr__res_xhigh_po W=0.69  L=4 mult=1 m=1
XM3 net3 net3 net2 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XM4 vd1 vd1 net3 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XM5 vd1 vd1 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XM6 vdd vd1 vssup vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XR4 vss vss vss sky130_fd_pr__res_xhigh_po W=0.69  L=4 mult=1 m=1
XR5 vss vss vss sky130_fd_pr__res_xhigh_po W=0.69  L=4 mult=1 m=1
.ends


* expanding   symbol:  Project/AR_BGR_with_Enable_line/schematic/fullldo/fullldoxc_v2_1.sym # of
*+ pins=7
** sym_path: /home/ahmedreda/Project/AR_BGR_with_Enable_line/schematic/fullldo/fullldoxc_v2_1.sym
** sch_path: /home/ahmedreda/Project/AR_BGR_with_Enable_line/schematic/fullldo/fullldoxc_v2_1.sch
.subckt fullldoxc_v2_1 trim[15] trim[14] trim[13] trim[12] trim[11] trim[10] trim[9] trim[8] trim[7]
+ trim[6] trim[5] trim[4] trim[3] trim[2] trim[1] trim[0] vss biasbgr vdd biasldo vg out
*.PININFO vss:B vdd:B biasldo:I out:O biasbgr:I trim[15:0]:I vg:O
XC2 gate vss sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=24 m=24
XC1 vref vss sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
x1 vdd vref vss biasbgr trim[15] trim[14] trim[13] trim[12] trim[11] trim[10] trim[9] trim[8]
+ trim[7] trim[6] trim[5] trim[4] trim[3] trim[2] trim[1] trim[0] gate bandgapxd
x2 vss vdd vg biasldo vref out ldoxc_1
.ends


* expanding   symbol:  Project/TG/tg1x.sym # of pins=4
** sym_path: /home/ahmedreda/Project/TG/tg1x.sym
** sch_path: /home/ahmedreda/Project/TG/tg1x.sch
.subckt tg1x vdd s vo vss
*.PININFO vdd:B vss:B s:I vo:O
XM1 sdash s vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM3 vdd sdash vo vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM4 sdash s vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM2 vdd s vo vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
.ends


* expanding   symbol:  Project/AR_BGR_with_Enable_line/schematic/bandgap_core/bandgapxd.sym # of
*+ pins=6
** sym_path: /home/ahmedreda/Project/AR_BGR_with_Enable_line/schematic/bandgap_core/bandgapxd.sym
** sch_path: /home/ahmedreda/Project/AR_BGR_with_Enable_line/schematic/bandgap_core/bandgapxd.sch
.subckt bandgapxd vdd vbg vss bias trim[15] trim[14] trim[13] trim[12] trim[11] trim[10] trim[9]
+ trim[8] trim[7] trim[6] trim[5] trim[4] trim[3] trim[2] trim[1] trim[0] gate
*.PININFO vbg:O bias:I trim[15:0]:I vdd:B vss:B gate:O
XM12 comp gate vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XM1 vbg gate vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XM2 vs2 vs2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XM6 vss vdd vs2 vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XC2 vs2 vss sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=4 m=4
XM3 vs1 vbg vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XM4 gate vs1 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
x2 vbg comp vp vn vss bg_res
x3 trimup veg trim[15] trim[14] trim[13] trim[12] trim[11] trim[10] trim[9] trim[8] trim[7] trim[6]
+ trim[5] trim[4] trim[3] trim[2] trim[1] trim[0] vss bg_trim
XQ1 vss vss vn sky130_fd_pr__pnp_05v5 W=0.68 L=0.68 m=1
XQ2 vss vss veg sky130_fd_pr__pnp_05v5 W=0.68 L=0.68 m=8
x7 vdd gate vp vn vss bias ota
XR2 trimup vp vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XM7 vdd vdd vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XR17 vss vss vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR18 vss vss vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR21 vss vss vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR23 vss vss vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XM5 vs1 vs2 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=1
.ends


* expanding   symbol:  Project/AR_BGR_with_Enable_line/schematic/ldo_core/ldoxc_1.sym # of pins=6
** sym_path: /home/ahmedreda/Project/AR_BGR_with_Enable_line/schematic/ldo_core/ldoxc_1.sym
** sch_path: /home/ahmedreda/Project/AR_BGR_with_Enable_line/schematic/ldo_core/ldoxc_1.sch
.subckt ldoxc_1 vss vdd vg bias vref out
*.PININFO out:O bias:I vss:B vdd:B vref:I vg:I
x3 vdd vg out pmosx
x1 vdd vg vref fbdiv bias vss otaldox
x2 out vss fbdiv vdx
XC4 vg out sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=20 m=20
XC5 out fbdiv sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=20 m=20
.ends


* expanding   symbol:  Project/AR_BGR/schematic/bandgap_core/bg_res.sym # of pins=5
** sym_path: /home/ahmedreda/Project/AR_BGR/schematic/bandgap_core/bg_res.sym
** sch_path: /home/ahmedreda/Project/AR_BGR/schematic/bandgap_core/bg_res.sch
.subckt bg_res b a d c vss
*.PININFO vss:B a:I b:I c:O d:O
XR21 net14 b vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR1 net15 net14 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR2 net16 net15 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR3 net17 net16 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR4 net18 net17 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR5 net6 net18 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR6 net8 net6 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR7 net10 net8 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR8 net12 net10 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR9 d net12 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR10 c net13 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR11 net13 net11 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR12 net7 net4 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR13 net9 net7 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR14 net11 net9 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR15 net4 net5 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR16 net5 net2 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR17 net2 net3 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR18 net3 net1 vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
XR19 net1 a vss sky130_fd_pr__res_xhigh_po W=0.69  L=13 mult=1 m=1
.ends


* expanding   symbol:  Project/AR_BGR/schematic/bandgap_core/bg_trim.sym # of pins=4
** sym_path: /home/ahmedreda/Project/AR_BGR/schematic/bandgap_core/bg_trim.sym
** sch_path: /home/ahmedreda/Project/AR_BGR/schematic/bandgap_core/bg_trim.sch
.subckt bg_trim top bot ctl[15] ctl[14] ctl[13] ctl[12] ctl[11] ctl[10] ctl[9] ctl[8] ctl[7] ctl[6]
+ ctl[5] ctl[4] ctl[3] ctl[2] ctl[1] ctl[0] vss
*.PININFO vss:B bot:B top:B ctl[15:0]:I
XM1 top ctl[15] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM2 net12 ctl[14] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM3 net11 ctl[13] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM4 net10 ctl[12] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM5 net9 ctl[11] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM6 net15 ctl[10] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM7 net14 ctl[9] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM8 net13 ctl[8] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM9 net6 ctl[5] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM10 net5 ctl[4] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM11 net7 ctl[6] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM12 net8 ctl[7] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM13 net3 ctl[2] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM14 net2 ctl[1] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM15 net1 ctl[0] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM16 net4 ctl[3] bot vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XR1 net12 top vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR2 net11 net12 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR3 net10 net11 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR4 net9 net10 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR5 net15 net9 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR6 net14 net15 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR7 net13 net14 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR8 net8 net13 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR9 net7 net8 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR10 net6 net7 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR11 net5 net6 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR12 net4 net5 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR13 net3 net4 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR14 net2 net3 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR15 net1 net2 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR16 bot net1 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
.ends


* expanding   symbol:  Project/AR_BGR/schematic/ota/ota.sym # of pins=6
** sym_path: /home/ahmedreda/Project/AR_BGR/schematic/ota/ota.sym
** sch_path: /home/ahmedreda/Project/AR_BGR/schematic/ota/ota.sch
.subckt ota vdd out inp inn vss bias
*.PININFO inn:I inp:I out:O bias:I vss:B vdd:B
XM12 vbp1 vbp1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM13 vbn2 vbp1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM14 bias1 bias1 vbp1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM1 outp inp diff vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=10
XM2 diff vbp1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=10
XM3 o1 vg vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM8 o2 vg vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM10 out bias1 o2 vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM11 vg bias1 o1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM19 vbn2 vbn2 vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM5 vg vbn2 outp vss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM9 outp vbn1 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=16
XM16 outn vbn1 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=16
XM7 out vbn2 outn vss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM6 vbn1 vbn1 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=4
XM15 outn inn diff vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=10
XM4 bias1 bias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=5 nf=1 m=2
XM17 bias bias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=5 nf=1 m=2
XM18 diff diff diff vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM20 vss vss vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=4
XM21 vss vss vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=4
XM22 vss vss vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=4
XM23 diff diff diff vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM24 vdd vdd vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM34 vbn1 vbn1 vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM33 bias1 bias1 bias1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM25 vg vg vg vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM26 out out out vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM27 out out out vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM28 vg vg vg vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=4
.ends


* expanding   symbol:  Project/AR_BGR/schematic/ldo_core/pmosx.sym # of pins=3
** sym_path: /home/ahmedreda/Project/AR_BGR/schematic/ldo_core/pmosx.sym
** sch_path: /home/ahmedreda/Project/AR_BGR/schematic/ldo_core/pmosx.sch
.subckt pmosx vdd vg vout
*.PININFO vout:O vdd:B vg:I
XM8 vout vg vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=44
XM1 vdd vdd vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=4
.ends


* expanding   symbol:  Project/AR_BGR/schematic/ldo_core/otaldox.sym # of pins=6
** sym_path: /home/ahmedreda/Project/AR_BGR/schematic/ldo_core/otaldox.sym
** sch_path: /home/ahmedreda/Project/AR_BGR/schematic/ldo_core/otaldox.sch
.subckt otaldox vdd otaout vref fbdiv bias vss
*.PININFO vref:I bias:I vss:B vdd:B fbdiv:I otaout:O
XM12 vbp1 vbp1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM13 vbn2 vbp1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM14 bias1 bias1 vbp1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM6 outp fbdiv diff vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=10
XM10 diff vbp1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=10
XM11 o1 vg vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM15 o2 vg vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM16 otaout bias1 o2 vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM17 vg bias1 o1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM19 vbn2 vbn2 vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM18 vg vbn2 outp vss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM20 outp vbn1 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=16
XM21 outn vbn1 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=16
XM22 otaout vbn2 outn vss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM23 vbn1 vbn1 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=4
XM24 outn vref diff vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=10
XM25 bias1 bias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=5 nf=1 m=2
XM26 bias bias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=5 nf=1 m=2
XM27 diff diff diff vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM28 vss vss vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=4
XM29 vss vss vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=4
XM30 vss vss vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=4
XM31 diff diff diff vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM32 vdd vdd vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM34 vbn1 vbn1 vbn1 vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM33 bias1 bias1 bias1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=4
XM35 vg vg vg vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM36 otaout otaout otaout vdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM37 otaout otaout otaout vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM38 vg vg vg vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=4
.ends


* expanding   symbol:  Project/AR_BGR/schematic/ldo_core/vdx.sym # of pins=3
** sym_path: /home/ahmedreda/Project/AR_BGR/schematic/ldo_core/vdx.sym
** sch_path: /home/ahmedreda/Project/AR_BGR/schematic/ldo_core/vdx.sch
.subckt vdx vout vss vb
*.PININFO vout:O vss:B vb:O
XR1 vb vout vss sky130_fd_pr__res_xhigh_po W=0.35 L=34 mult=1 m=1
XR2 vss vb vss sky130_fd_pr__res_xhigh_po W=0.35 L=34 mult=1 m=1
XR3 vss vss vss sky130_fd_pr__res_xhigh_po W=0.35 L=8.5 mult=1 m=1
XR4 vss vss vss sky130_fd_pr__res_xhigh_po W=0.35 L=8.5 mult=1 m=1
XR5 vb vout vss sky130_fd_pr__res_xhigh_po W=0.35 L=34 mult=1 m=1
.ends

.end